// Copyright(C) 2020-2022 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by MIT and ISC licenses (mapbox).
// Both files are distributed with this software package.
module main

import earcut

fn main() {
	flat_dude := earcut.flatten(dude)
	vertices := flat_dude.vertices
	holes := flat_dude.holes
	indicies := earcut.earcut(vertices, holes, 2)
	println(earcut.deviation(vertices, holes, 2, indicies))
}

const dude = [
	[
		[f32(280.35714), 648.79075],
		[f32(286.78571), 662.8979],
		[f32(263.28607), 661.17871],
		[f32(262.31092), 671.41548],
		[f32(250.53571), 677.00504],
		[f32(250.53571), 683.43361],
		[f32(256.42857), 685.21933],
		[f32(297.14286), 669.50504],
		[f32(289.28571), 649.50504],
		[f32(285), 631.6479],
		[f32(285), 608.79075],
		[f32(292.85714), 585.21932],
		[f32(306.42857), 563.79075],
		[f32(323.57143), 548.79075],
		[f32(339.28571), 545.21932],
		[f32(357.85714), 547.36218],
		[f32(375), 550.21932],
		[f32(391.42857), 568.07647],
		[f32(404.28571), 588.79075],
		[f32(413.57143), 612.36218],
		[f32(417.14286), 628.07647],
		[f32(438.57143), 619.1479],
		[f32(438.03572), 618.96932],
		[f32(437.5), 609.50504],
		[f32(426.96429), 609.86218],
		[f32(424.64286), 615.57647],
		[f32(419.82143), 615.04075],
		[f32(420.35714), 605.04075],
		[f32(428.39286), 598.43361],
		[f32(437.85714), 599.68361],
		[f32(443.57143), 613.79075],
		[f32(450.71429), 610.21933],
		[f32(431.42857), 575.21932],
		[f32(405.71429), 550.21932],
		[f32(372.85714), 534.50504],
		[f32(349.28571), 531.6479],
		[f32(346.42857), 521.6479],
		[f32(346.42857), 511.6479],
		[f32(350.71429), 496.6479],
		[f32(367.85714), 476.6479],
		[f32(377.14286), 460.93361],
		[f32(385.71429), 445.21932],
		[f32(388.57143), 404.50504],
		[f32(360), 352.36218],
		[f32(337.14286), 325.93361],
		[f32(330.71429), 334.50504],
		[f32(347.14286), 354.50504],
		[f32(337.85714), 370.21932],
		[f32(333.57143), 359.50504],
		[f32(319.28571), 353.07647],
		[f32(312.85714), 366.6479],
		[f32(350.71429), 387.36218],
		[f32(368.57143), 408.07647],
		[f32(375.71429), 431.6479],
		[f32(372.14286), 454.50504],
		[f32(366.42857), 462.36218],
		[f32(352.85714), 462.36218],
		[f32(336.42857), 456.6479],
		[f32(332.85714), 438.79075],
		[f32(338.57143), 423.79075],
		[f32(338.57143), 411.6479],
		[f32(327.85714), 405.93361],
		[f32(320.71429), 407.36218],
		[f32(315.71429), 423.07647],
		[f32(314.28571), 440.21932],
		[f32(325), 447.71932],
		[f32(324.82143), 460.93361],
		[f32(317.85714), 470.57647],
		[f32(304.28571), 483.79075],
		[f32(287.14286), 491.29075],
		[f32(263.03571), 498.61218],
		[f32(251.60714), 503.07647],
		[f32(251.25), 533.61218],
		[f32(260.71429), 533.61218],
		[f32(272.85714), 528.43361],
		[f32(286.07143), 518.61218],
		[f32(297.32143), 508.25504],
		[f32(297.85714), 507.36218],
		[f32(298.39286), 506.46932],
		[f32(307.14286), 496.6479],
		[f32(312.67857), 491.6479],
		[f32(317.32143), 503.07647],
		[f32(322.5), 514.1479],
		[f32(325.53571), 521.11218],
		[f32(327.14286), 525.75504],
		[f32(326.96429), 535.04075],
		[f32(311.78571), 540.04075],
		[f32(291.07143), 552.71932],
		[f32(274.82143), 568.43361],
		[f32(259.10714), 592.8979],
		[f32(254.28571), 604.50504],
		[f32(251.07143), 621.11218],
		[f32(250.53571), 649.1479],
		[f32(268.1955), 654.36208],
	],
	[
		[f32(325), 437],
		[f32(320), 423],
		[f32(329), 413],
		[f32(332), 423],
	],
	[
		[f32(320.72342), 480],
		[f32(338.90617), 465.96863],
		[f32(347.99754), 480.61584],
		[f32(329.8148), 510.41534],
		[f32(339.91632), 480.11077],
		[f32(334.86556), 478.09046],
	],
]
